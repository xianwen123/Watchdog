`ifndef RKV_WATCHDOG_ELEMENT_SEQUENCES_SVH
`define RKV_WATCHDOG_ELEMENT_SEQUENCES_SVH


`include "rkv_watchdog_base_element_sequence.sv"
`include "rkv_watchdog_reg_enable_intr.sv"
`include "rkv_watchdog_reg_disable_intr.sv"
`include "rkv_watchdog_reg_enable_reset.sv"
`include "rkv_watchdog_reg_loadcount.sv"
`include "rkv_watchdog_reg_intr_wait_clear.sv"


`endif // RKV_WATCHDOG_ELEMENT_SEQUENCES_SVH
