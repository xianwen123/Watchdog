`ifndef RKV_WATCHDOG_REG_SVH
`define RKV_WATCHDOG_REG_SVH

`include "rkv_watchdog_reg.sv"

`endif // RKV_WATCHDOG_REG_SVH
